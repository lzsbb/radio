domain gateway broadcast
