nameserver 10.0.0.138
search gateway
